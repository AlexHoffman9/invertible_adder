// Alex Hoffman, McGill University
// outputs a stochastic "p-bit:" a biased random bit depending on the outputs of its neighbors
module pbit(clk, reset, p_in, I_0, update_control, clamp_control, p_out);
parameter SEED = 32'h98390184,      // SEED for prng
N_NEIGHBORS = 4,                    // number of pbit connections
WEIGHT_PRECISION = 6,               // bit precision of weights, tanh input
H = 6'd1,                           // constant offset for this pbit
W = {6'd1, 6'd1, 6'd1, 6'd1},       // weights for this pbit in s[3][2] format -8 to 7.75 range for tanh input
WIDTH = 8;

input clk, reset, update_control;   // clk, reset, update_control==1 allows pbit to update its output, otherwise it holds
input[N_NEIGHBORS-1:0] p_in;        // input p bits
input [3:0] I_0;                    // unsigned scaling. fixed point [2][2]
input [1:0] clamp_control;          // msb = clamp enable, lsb = clamped value
output reg p_out;                   // output bit

// local vars to connect modules
wire[5:0] I_i;                      // output of MAC, input to activation function
wire[WIDTH-1:0] activation;              // output of activation function
wire[WIDTH-1:0] sum;                     // sum of prng and activation output. The output is drawn from the sign of this sum
wire[WIDTH-1:0] prng_out;                // pseudo random number generated by lfsr

// prng
// prng_32 prng(clk, reset, SEED, prng_out);
prng_8 prng(clk,reset,SEED,prng_out);

// MAC. Outputs weighted sum of input pbits, thresholded to 6 bits
mac #(N_NEIGHBORS, WEIGHT_PRECISION, H, W) mac_pbit(p_in, I_0, I_i);

// tanh. inputs: I_i (MAC output), outputs: activation
// tanh tan(I_i, activation); // LUT TANH
fast_tanh #(WIDTH) tan(I_i, activation);

// combinational logic for sum of random number and activation output
assign sum = prng_out+activation; 

// sequential logic for updating output bit
always@(posedge clk) begin
    if (clamp_control[1]) begin // if pbit output should be clamped to a value (this pbit acts as input to boltzmann machine)
        p_out <= clamp_control[0];
    end else if (reset) begin
        p_out <= SEED[WIDTH-1];      // random reset bit
    end else begin 
        if (update_control) begin // update pbit when high
            p_out <= ~(prng_out[WIDTH-1]&activation[WIDTH-1] || ((prng_out[WIDTH-1]^activation[WIDTH-1])&sum[WIDTH-1]));  // if sum is negative (operands are pos or operands are pos,neg and num to pos)
        end else begin // pbit should not be updated
            p_out <= p_out;
        end
    end
end
endmodule


`timescale 1ns/1ps
module pbit_testbench();
localparam N_NEIGHBORS = 4, WEIGHT_PRECISION = 6, SEED = 32'h48390184, H = 6'd0, W = {6'd3, 6'd2, -6'd1, -6'd1}, WIDTH = 32; 
reg clk, reset;
reg[N_NEIGHBORS-1:0] p_in;    // input p bits
reg [3:0] I_0;
wire p_out;                   // output bit
reg update_control;
reg [1:0] clamp_control; 

pbit #(SEED, N_NEIGHBORS, WEIGHT_PRECISION, H, W, WIDTH) dut(clk, reset, p_in, I_0, update_control, clamp_control, p_out);

parameter CLOCK_PERIOD = 20;
	initial // Clock setUp
	begin
		clk = 0; 
		forever #(CLOCK_PERIOD/2) clk <= ~clk;
	end

integer i; integer sum = 0; integer steps = 100;
initial 
begin
    reset <= 1; I_0 <= 4'd4; p_in <= 4'b0000; clamp_control <= 2'b00; update_control <= 1'b1;
    #CLOCK_PERIOD; reset <= 0;#CLOCK_PERIOD; reset <= 1;#CLOCK_PERIOD; reset <= 0;
    for (i = 0; i < steps; i = i + 1) begin 
        #CLOCK_PERIOD;
        p_in <= p_in + 1;
    end


    // #CLOCK_PERIOD; #CLOCK_PERIOD; #CLOCK_PERIOD; #CLOCK_PERIOD; clamp_control <= 2'b10;
    // #CLOCK_PERIOD; #CLOCK_PERIOD; #CLOCK_PERIOD; #CLOCK_PERIOD; clamp_control <= 2'b11;
    // #CLOCK_PERIOD; #CLOCK_PERIOD; #CLOCK_PERIOD; #CLOCK_PERIOD; clamp_control <= 2'b01;
    // #CLOCK_PERIOD; #CLOCK_PERIOD; #CLOCK_PERIOD; #CLOCK_PERIOD; clamp_control <= 2'b01;
    // #CLOCK_PERIOD; #CLOCK_PERIOD; #CLOCK_PERIOD; #CLOCK_PERIOD; update_control <= 1'b0;
    for (i = 0; i < 16; i = i + 1) begin 
        #CLOCK_PERIOD;
        sum = sum + 2*p_out - 1;
    end
    $display("input weights = %b, average value = %f after %d bits", p_in, sum*1.0/steps, steps);
    // $display("expected average value for tanh input %d is %f", 1, 0.76);

    // p_in <= 4'b1110;sum=0;
    // for (i = 0; i < steps; i = i + 1) begin 
    //     #CLOCK_PERIOD;
    //     sum = sum + 2*p_out - 1;
    // end
    // $display("input weights = %b, average value = %f after %d bits", p_in, sum*1.0/steps, steps);
    // p_in <= 4'b1100; sum=0;
    // for (i = 0; i < steps; i = i + 1) begin 
    //     #CLOCK_PERIOD;
    //     sum = sum + 2*p_out - 1;
    // end
    // $display("input weights = %b, average value = %f after %d bits", p_in, sum*1.0/steps, steps);
    // p_in <= 4'b1000;sum=0;
    // for (i = 0; i < steps; i = i + 1) begin 
    //     #CLOCK_PERIOD;
    //     sum = sum + 2*p_out - 1;
    // end
    // $display("input weights = %b, average value = %f after %d bits", p_in, sum*1.0/steps, steps);
    //  p_in <= 4'b0000;sum=0;
    // for (i = 0; i < steps; i = i + 1) begin 
    //     #CLOCK_PERIOD;
    //     sum = sum + 2*p_out - 1;
    // end
    // $display("input weights = %b, average value = %f after %d bits", p_in, sum*1.0/steps, steps);
    $stop;
end
endmodule