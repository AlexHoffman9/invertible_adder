// Alex Hoffman, McGill University
// tanh function implemented with lookup table
// 6 bit address and 32 bit output s[31] fixed point format
module tanh(in, out);
input[5:0] in;  // 6 bits 2's complement fixed point. s[3][2] format
output reg[31:0] out; // 32 bit 2's comp output -1 to (almost) 1 range

always @(*)
begin
    case (in)
        -6'd32: out = -32'd2147483164;
        -6'd31: out = -32'd2147482851;
        -6'd30: out = -32'd2147482334;
        -6'd29: out = -32'd2147481481;
        -6'd28: out = -32'd2147480076;
        -6'd27: out = -32'd2147477759;
        -6'd26: out = -32'd2147473939;
        -6'd25: out = -32'd2147467642;
        -6'd24: out = -32'd2147457258;
        -6'd23: out = -32'd2147440140;
        -6'd22: out = -32'd2147411915;
        -6'd21: out = -32'd2147365383;
        -6'd20: out = -32'd2147288665;
        -6'd19: out = -32'd2147162185;
        -6'd18: out = -32'd2146953672;
        -6'd17: out = -32'd2146609935;
        -6'd16: out = -32'd2146043330;
        -6'd15: out = -32'd2145109481;
        -6'd14: out = -32'd2143570712;
        -6'd13: out = -32'd2141036119;
        -6'd12: out = -32'd2136863812;
        -6'd11: out = -32'd2130002539;
        -6'd10: out = -32'd2118738072;
        -6'd9: out = -32'd2100295088;
        -6'd8: out = -32'd2070233464;
        -6'd7: out = -32'd2021588575;
        -6'd6: out = -32'd1943791073;
        -6'd5: out = -32'd1821675245;
        -6'd4: out = -32'd1635510996;
        -6'd3: out = -32'd1363971989;
        -6'd2: out = -32'd992389038;
        -6'd1: out = -32'd525958822;
        6'd0: out = 32'd0;
        6'd1: out = 32'd525958822;
        6'd2: out = 32'd992389038;
        6'd3: out = 32'd1363971989;
        6'd4: out = 32'd1635510996;
        6'd5: out = 32'd1821675245;
        6'd6: out = 32'd1943791073;
        6'd7: out = 32'd2021588575;
        6'd8: out = 32'd2070233464;
        6'd9: out = 32'd2100295088;
        6'd10: out = 32'd2118738072;
        6'd11: out = 32'd2130002539;
        6'd12: out = 32'd2136863812;
        6'd13: out = 32'd2141036119;
        6'd14: out = 32'd2143570712;
        6'd15: out = 32'd2145109481;
        6'd16: out = 32'd2146043330;
        6'd17: out = 32'd2146609935;
        6'd18: out = 32'd2146953672;
        6'd19: out = 32'd2147162185;
        6'd20: out = 32'd2147288665;
        6'd21: out = 32'd2147365383;
        6'd22: out = 32'd2147411915;
        6'd23: out = 32'd2147440140;
        6'd24: out = 32'd2147457258;
        6'd25: out = 32'd2147467642;
        6'd26: out = 32'd2147473939;
        6'd27: out = 32'd2147477759;
        6'd28: out = 32'd2147480076;
        6'd29: out = 32'd2147481481;
        6'd30: out = 32'd2147482334;
        6'd31: out = 32'd2147482851;
        default: out <= 32'd1;
    endcase
end
endmodule