// Alex Hoffman, McGill University
// tanh function implemented with lookup table
// 6 bit address and 32 bit output s[31] fixed point format
module tanh(in, out);
input[5:0] in;  // 6 bits 2's complement fixed point. s[3][2] format
output reg[31:0] out; // 32 bit 2's comp output -1 to (almost) 1 range

always @(*)
begin
    case (in)
        -6'd32: out = -32'd1073741582;
        -6'd31: out = -32'd1073741425;
        -6'd30: out = -32'd1073741167;
        -6'd29: out = -32'd1073740740;
        -6'd28: out = -32'd1073740038;
        -6'd27: out = -32'd1073738879;
        -6'd26: out = -32'd1073736969;
        -6'd25: out = -32'd1073733821;
        -6'd24: out = -32'd1073728629;
        -6'd23: out = -32'd1073720070;
        -6'd22: out = -32'd1073705957;
        -6'd21: out = -32'd1073682691;
        -6'd20: out = -32'd1073644332;
        -6'd19: out = -32'd1073581092;
        -6'd18: out = -32'd1073476836;
        -6'd17: out = -32'd1073304967;
        -6'd16: out = -32'd1073021665;
        -6'd15: out = -32'd1072554740;
        -6'd14: out = -32'd1071785356;
        -6'd13: out = -32'd1070518059;
        -6'd12: out = -32'd1068431906;
        -6'd11: out = -32'd1065001269;
        -6'd10: out = -32'd1059369036;
        -6'd9: out = -32'd1050147544;
        -6'd8: out = -32'd1035116732;
        -6'd7: out = -32'd1010794287;
        -6'd6: out = -32'd971895536;
        -6'd5: out = -32'd910837622;
        -6'd4: out = -32'd817755498;
        -6'd3: out = -32'd681985994;
        -6'd2: out = -32'd496194519;
        -6'd1: out = -32'd262979411;
        6'd0: out = 32'd0;
        6'd1: out = 32'd262979411;
        6'd2: out = 32'd496194519;
        6'd3: out = 32'd681985994;
        6'd4: out = 32'd817755498;
        6'd5: out = 32'd910837622;
        6'd6: out = 32'd971895536;
        6'd7: out = 32'd1010794287;
        6'd8: out = 32'd1035116732;
        6'd9: out = 32'd1050147544;
        6'd10: out = 32'd1059369036;
        6'd11: out = 32'd1065001269;
        6'd12: out = 32'd1068431906;
        6'd13: out = 32'd1070518059;
        6'd14: out = 32'd1071785356;
        6'd15: out = 32'd1072554740;
        6'd16: out = 32'd1073021665;
        6'd17: out = 32'd1073304967;
        6'd18: out = 32'd1073476836;
        6'd19: out = 32'd1073581092;
        6'd20: out = 32'd1073644332;
        6'd21: out = 32'd1073682691;
        6'd22: out = 32'd1073705957;
        6'd23: out = 32'd1073720070;
        6'd24: out = 32'd1073728629;
        6'd25: out = 32'd1073733821;
        6'd26: out = 32'd1073736969;
        6'd27: out = 32'd1073738879;
        6'd28: out = 32'd1073740038;
        6'd29: out = 32'd1073740740;
        6'd30: out = 32'd1073741167;
        6'd31: out = 32'd1073741425;
        default: out <= 32'd1;
    endcase
end
endmodule